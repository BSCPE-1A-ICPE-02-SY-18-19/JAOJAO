CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
11
7 Ground~
168 854 28 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5130 0 0
2
43530.3 0
0
2 +V
167 175 158 0 1 3
0 16
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
391 0 0
2
43530.3 0
0
9 2-In AND~
219 483 97 0 3 22
0 15 11 14
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3124 0 0
2
43530.3 0
0
9 2-In AND~
219 356 96 0 3 22
0 13 12 15
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3421 0 0
2
43530.3 0
0
9 CC 7-Seg~
183 860 114 0 17 19
10 3 4 5 6 7 8 9 18 2
0 0 0 1 1 0 1 2
0
0 0 21088 0
6 BLUECC
13 -41 55 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
8157 0 0
2
43530.3 0
0
6 74LS48
188 694 177 0 14 29
0 10 11 12 13 19 20 9 8 7
6 5 4 3 21
0
0 0 4848 0
6 74LS48
-21 -60 21 -52
2 U3
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 0 0 0 0
1 U
5572 0 0
2
43530.3 0
0
6 74112~
219 528 258 0 7 32
0 16 14 17 14 16 10 22
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
8901 0 0
2
43530.3 0
0
6 74112~
219 415 259 0 7 32
0 16 15 17 15 16 23 11
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
7361 0 0
2
43530.3 0
0
6 74112~
219 288 260 0 7 32
0 16 13 17 13 16 24 12
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U1B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
4747 0 0
2
43530.3 0
0
6 74112~
219 175 261 0 7 32
0 16 25 17 26 16 27 13
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U1A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
972 0 0
2
43530.3 0
0
7 Pulser~
4 55 284 0 10 12
0 28 29 30 17 0 0 5 5 2
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
3472 0 0
2
43530.3 0
0
36
1 9 2 0 0 12416 0 1 5 0 0 6
854 22
854 18
868 18
868 64
860 64
860 72
13 1 3 0 0 4224 0 6 5 0 0 3
726 195
839 195
839 150
12 2 4 0 0 4224 0 6 5 0 0 3
726 186
845 186
845 150
11 3 5 0 0 4224 0 6 5 0 0 3
726 177
851 177
851 150
10 4 6 0 0 4224 0 6 5 0 0 3
726 168
857 168
857 150
9 5 7 0 0 4224 0 6 5 0 0 3
726 159
863 159
863 150
8 6 8 0 0 4224 0 6 5 0 0 5
726 150
825 150
825 163
869 163
869 150
7 7 9 0 0 4224 0 6 5 0 0 5
726 141
830 141
830 158
875 158
875 150
6 1 10 0 0 8320 0 7 6 0 0 4
558 240
654 240
654 141
662 141
0 2 11 0 0 4224 0 0 6 15 0 2
451 150
662 150
0 3 12 0 0 4224 0 0 6 19 0 2
324 159
662 159
0 4 13 0 0 8320 0 0 6 22 0 3
248 225
248 168
662 168
0 2 14 0 0 12288 0 0 7 14 0 6
493 225
562 225
562 185
490 185
490 222
504 222
3 4 14 0 0 8320 0 3 7 0 0 6
504 97
508 97
508 191
493 191
493 240
504 240
7 2 11 0 0 0 0 8 3 0 0 4
439 223
451 223
451 106
459 106
0 2 15 0 0 8192 0 0 8 18 0 3
381 223
381 223
391 223
0 1 15 0 0 4096 0 0 3 18 0 4
381 98
451 98
451 88
459 88
4 3 15 0 0 8320 0 8 4 0 0 4
391 241
381 241
381 96
377 96
7 2 12 0 0 0 0 9 4 0 0 4
312 224
324 224
324 105
332 105
0 1 13 0 0 0 0 0 4 21 0 4
258 196
254 196
254 87
332 87
0 4 13 0 0 0 0 0 9 22 0 5
258 224
258 193
240 193
240 242
264 242
7 2 13 0 0 0 0 10 9 0 0 4
199 225
250 225
250 224
264 224
0 0 16 0 0 4096 0 0 0 28 32 2
466 176
466 278
0 0 16 0 0 0 0 0 0 28 32 2
348 176
348 278
0 0 16 0 0 0 0 0 0 28 32 2
234 176
234 278
0 1 16 0 0 0 0 0 8 28 0 4
416 176
416 188
415 188
415 196
0 1 16 0 0 0 0 0 9 28 0 2
288 176
288 197
0 1 16 0 0 4224 0 0 7 29 0 3
175 176
528 176
528 195
1 1 16 0 0 0 0 2 10 0 0 2
175 167
175 198
5 0 16 0 0 0 0 8 0 0 32 3
415 271
415 278
416 278
5 0 16 0 0 0 0 9 0 0 32 3
288 272
288 278
289 278
5 5 16 0 0 0 0 10 7 0 0 4
175 273
175 278
528 278
528 270
0 3 17 0 0 4096 0 0 8 36 0 3
359 284
359 232
385 232
0 3 17 0 0 0 0 0 9 36 0 3
244 284
244 233
258 233
0 3 17 0 0 0 0 0 10 36 0 3
119 284
119 234
145 234
4 3 17 0 0 4224 0 11 7 0 0 4
85 284
490 284
490 231
498 231
1
-16 0 0 0 700 0 0 0 0 3 2 1 66
11 Kristen ITC
0 0 0 20
182 313 440 348
193 321 428 344
20 JAOJAO, CARL JOHN E.
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
